package cmd_bits;

	// command bit description
	localparam b_tx = 0, b_op_1 = 1, b_op_2 = 2, b_subres = 4, b_addres = 5, b_subop = 6, b_addop = 7;

endpackage